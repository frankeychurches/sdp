module hex7seg (input )