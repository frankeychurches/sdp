module adder_4b (sum