module luces_fsm (
    clk, reset, enable, leds
);


input clk, reset, enable;
output [7:0] leds;

parameter  = ;
    
endmodule